//--------------------------------------------------------------------------------------------
// Module: Hvl top module
//--------------------------------------------------------------------------------------------
module hvl_top;

  //-------------------------------------------------------
  // Package : Importing Uvm Pakckage and Test Package
  //-------------------------------------------------------
  import test_pkg::*;
  import uvm_pkg::*;

  //-------------------------------------------------------
  // Declaring UART Interface
  //-------------------------------------------------------
  //uart_if vif();

  //-------------------------------------------------------
  // run_test for simulation
  //-------------------------------------------------------
  initial begin
    //-------------------------------------------------------
    // Setting UART Interface
    //-------------------------------------------------------
    //uvm_config_db #(virtual uart_if)::set(null,"*","vif",vif); 
    run_test("base_test");
  end

endmodule : hvl_top
